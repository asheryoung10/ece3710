module seven_seg_decoder (
    input  wire [3:0] bin,   // 4-bit binary input
    output reg  [6:0] hex    // 7-seg output (active LOW)
);

    always @(*) begin
        case (bin)
            4'h0: hex = 7'b1000000; // 0
            4'h1: hex = 7'b1111001; // 1
            4'h2: hex = 7'b0100100; // 2
            4'h3: hex = 7'b0110000; // 3
            4'h4: hex = 7'b0011001; // 4
            4'h5: hex = 7'b0010010; // 5
            4'h6: hex = 7'b0000010; // 6
            4'h7: hex = 7'b1111000; // 7
            4'h8: hex = 7'b0000000; // 8
            4'h9: hex = 7'b0010000; // 9
            4'hA: hex = 7'b0001000; // A
            4'hB: hex = 7'b0000011; // b
            4'hC: hex = 7'b1000110; // C
            4'hD: hex = 7'b0100001; // d
            4'hE: hex = 7'b0000110; // E
            4'hF: hex = 7'b0001110; // F
            default: hex = 7'b1111111; // all OFF
        endcase
    end

endmodule
